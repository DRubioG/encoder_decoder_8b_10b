library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity decoder_8b_10b is
    Port (  
        clk : in std_logic;
        rst_n : in std_logic;
        data_in_p : in std_logic_vector(9 downto 0);
        data_in_n : in std_logic_vector(9 downto 0); -- diff positive
        data_out : out std_logic_vector(7 downto 0)  -- diff negative
    );
end decoder_8b_10b;

architecture arch_decoder_8b_10b of decoder_8b_10b is

signal data_out_aux, data_out_aux_2 : std_logic_vector(7 downto 0);

begin
    process (clk, rst_n, data_in_p)
    begin
        if rst_n = '0' then
            data_out_aux <= (others=>'0');
        elsif rising_edge(clk) then
            case data_in_p is
                when "0110001011" =>  -- D0.0
                    data_out_aux <= "00000000";
                when "1000101011" =>  -- D1.0
                    data_out_aux <= "00000001";
                when "0100101011" =>  -- D2.0
                    data_out_aux <= "00000010";
                when "1100010100" =>  -- D3.0
                    data_out_aux <= "00000011";
                when "0010101011" =>  -- D4.0
                    data_out_aux <= "00000100";
                when "1010010100" =>  -- D5.0
                    data_out_aux <= "00000101";
                when "0110010100" =>  -- D6.0
                    data_out_aux <= "00000110";
                when "0001110100" =>  -- D7.0
                    data_out_aux <= "00000111";
                when "0001101011" =>  -- D8.0
                    data_out_aux <= "00001000";
                when "1001010100" =>  -- D9.0
                    data_out_aux <= "00001001";
                when "0101010100" =>  -- D10.0
                    data_out_aux <= "00001010";
                when "1101000100" =>  -- D11.0
                    data_out_aux <= "00001011";
                when "0011010100" =>  -- D12.0
                    data_out_aux <= "00001100";
                when "1011000100" =>  -- D13.0
                    data_out_aux <= "00001101";
                when "0111000100" =>  -- D14.0
                    data_out_aux <= "00001110";
                when "1010001011" =>  -- D15.0
                    data_out_aux <= "00001111";
                when "1001001011" =>  -- D16.0
                    data_out_aux <= "00010000";
                when "1000110100" =>  -- D17.0
                    data_out_aux <= "00010001";
                when "0100110100" =>  -- D18.0
                    data_out_aux <= "00010010";
                when "1100100100" =>  -- D19.0
                    data_out_aux <= "00010011";
                when "0010110100" =>  -- D20.0
                    data_out_aux <= "00010100";
                when "1010100100" =>  -- D21.0
                    data_out_aux <= "00010101";
                when "0110100100" =>  -- D22.0
                    data_out_aux <= "00010110";
                when "0001011011" =>  -- D23.0
                    data_out_aux <= "00010111";
                when "0011001011" =>  -- D24.0
                    data_out_aux <= "00011000";
                when "1001100100" =>  -- D25.0
                    data_out_aux <= "00011001";
                when "0101100100" =>  -- D26.0
                    data_out_aux <= "00011010";
                when "0010011011" =>  -- D27.0
                    data_out_aux <= "00011011";
                when "0011100100" =>  -- D28.0
                    data_out_aux <= "00011100";
                when "0100011011" =>  -- D29.0
                    data_out_aux <= "00011101";
                when "1000011011" =>  -- D30.0
                    data_out_aux <= "00011110";
                when "0101001011" =>  -- D31.0
                    data_out_aux <= "00011111";
                when "0110001001" =>  -- D0.1
                    data_out_aux <= "00100000";
                when "1000101001" =>  -- D1.1
                    data_out_aux <= "00100001";
                when "0100101001" =>  -- D2.1
                    data_out_aux <= "00100010";
                when "1100011001" =>  -- D3.1
                    data_out_aux <= "00100011";
                when "0010101001" =>  -- D4.1
                    data_out_aux <= "00100100";
                when "1010011001" =>  -- D5.1
                    data_out_aux <= "00100101";
                when "0110011001" =>  -- D6.1
                    data_out_aux <= "00100110";
                when "0001111001" =>  -- D7.1
                    data_out_aux <= "00100111";
                when "0001101001" =>  -- D8.1
                    data_out_aux <= "00101000";
                when "1001011001" =>  -- D9.1
                    data_out_aux <= "00101001";
                when "0101011001" =>  -- D10.1
                    data_out_aux <= "00101010";
                when "1101001001" =>  -- D11.1
                    data_out_aux <= "00101011";
                when "0011011001" =>  -- D12.1
                    data_out_aux <= "00101100";
                when "1011001001" =>  -- D13.1
                    data_out_aux <= "00101101";
                when "0111001001" =>  -- D14.1
                    data_out_aux <= "00101110";
                when "1010001001" =>  -- D15.1
                    data_out_aux <= "00101111";
                when "1001001001" =>  -- D16.1
                    data_out_aux <= "00110000";
                when "1000111001" =>  -- D17.1
                    data_out_aux <= "00110001";
                when "0100111001" =>  -- D18.1
                    data_out_aux <= "00110010";
                when "1100101001" =>  -- D19.1
                    data_out_aux <= "00110011";
                when "0010111001" =>  -- D20.1
                    data_out_aux <= "00110100";
                when "1010101001" =>  -- D21.1
                    data_out_aux <= "00110101";
                when "0110101001" =>  -- D22.1
                    data_out_aux <= "00110110";
                when "0001011001" =>  -- D23.1
                    data_out_aux <= "00110111";
                when "0011001001" =>  -- D24.1
                    data_out_aux <= "00111000";
                when "1001101001" =>  -- D25.1
                    data_out_aux <= "00111001";
                when "0101101001" =>  -- D26.1
                    data_out_aux <= "00111010";
                when "0010011001" =>  -- D27.1
                    data_out_aux <= "00111011";
                when "0011101001" =>  -- D28.1
                    data_out_aux <= "00111100";
                when "0100011001" =>  -- D29.1
                    data_out_aux <= "00111101";
                when "1000011001" =>  -- D30.1
                    data_out_aux <= "00111110";
                when "0101001001" =>  -- D31.1
                    data_out_aux <= "00111111";
                when "0110000101" =>  -- D0.2
                    data_out_aux <= "01000000";
                when "1000100101" =>  -- D1.2
                    data_out_aux <= "01000001";
                when "0100100101" =>  -- D2.2
                    data_out_aux <= "01000010";
                when "1100010101" =>  -- D3.2
                    data_out_aux <= "01000011";
                when "0010100101" =>  -- D4.2
                    data_out_aux <= "01000100";
                when "1010010101" =>  -- D5.2
                    data_out_aux <= "01000101";
                when "0110010101" =>  -- D6.2
                    data_out_aux <= "01000110";
                when "0001110101" =>  -- D7.2
                    data_out_aux <= "01000111";
                when "0001100101" =>  -- D8.2
                    data_out_aux <= "01001000";
                when "1001010101" =>  -- D9.2
                    data_out_aux <= "01001001";
                when "0101010101" =>  -- D10.2
                    data_out_aux <= "01001010";
                when "1101000101" =>  -- D11.2
                    data_out_aux <= "01001011";
                when "0011010101" =>  -- D12.2
                    data_out_aux <= "01001100";
                when "1011000101" =>  -- D13.2
                    data_out_aux <= "01001101";
                when "0111000101" =>  -- D14.2
                    data_out_aux <= "01001110";
                when "1010000101" =>  -- D15.2
                    data_out_aux <= "01001111";
                when "1001000101" =>  -- D16.2
                    data_out_aux <= "01010000";
                when "1000110101" =>  -- D17.2
                    data_out_aux <= "01010001";
                when "0100110101" =>  -- D18.2
                    data_out_aux <= "01010010";
                when "1100100101" =>  -- D19.2
                    data_out_aux <= "01010011";
                when "0010110101" =>  -- D20.2
                    data_out_aux <= "01010100";
                when "1010100101" =>  -- D21.2
                    data_out_aux <= "01010101";
                when "0110100101" =>  -- D22.2
                    data_out_aux <= "01010110";
                when "0001010101" =>  -- D23.2
                    data_out_aux <= "01010111";
                when "0011000101" =>  -- D24.2
                    data_out_aux <= "01011000";
                when "1001100101" =>  -- D25.2
                    data_out_aux <= "01011001";
                when "0101100101" =>  -- D26.2
                    data_out_aux <= "01011010";
                when "0010010101" =>  -- D27.2
                    data_out_aux <= "01011011";
                when "0011100101" =>  -- D28.2
                    data_out_aux <= "01011100";
                when "0100010101" =>  -- D29.2
                    data_out_aux <= "01011101";
                when "1000010101" =>  -- D30.2
                    data_out_aux <= "01011110";
                when "0101000101" =>  -- D31.2
                    data_out_aux <= "01011111";
                when "0110001100" =>  -- D0.3
                    data_out_aux <= "01100000";
                when "1000101100" =>  -- D1.3
                    data_out_aux <= "01100001";
                when "0100101100" =>  -- D2.3
                    data_out_aux <= "01100010";
                when "1100010011" =>  -- D3.3
                    data_out_aux <= "01100011";
                when "0010101100" =>  -- D4.3
                    data_out_aux <= "01100100";
                when "1010010011" =>  -- D5.3
                    data_out_aux <= "01100101";
                when "0110010011" =>  -- D6.3
                    data_out_aux <= "01100110";
                when "0001110011" =>  -- D7.3
                    data_out_aux <= "01100111";
                when "0001101100" =>  -- D8.3
                    data_out_aux <= "01101000";
                when "1001010011" =>  -- D9.3
                    data_out_aux <= "01101001";
                when "0101010011" =>  -- D10.3
                    data_out_aux <= "01101010";
                when "1101000011" =>  -- D11.3
                    data_out_aux <= "01101011";
                when "0011010011" =>  -- D12.3
                    data_out_aux <= "01101100";
                when "1011000011" =>  -- D13.3
                    data_out_aux <= "01101101";
                when "0111000011" =>  -- D14.3
                    data_out_aux <= "01101110";
                when "1010001100" =>  -- D15.3
                    data_out_aux <= "01101111";
                when "1001001100" =>  -- D16.3
                    data_out_aux <= "01110000";
                when "1000110011" =>  -- D17.3
                    data_out_aux <= "01110001";
                when "0100110011" =>  -- D18.3
                    data_out_aux <= "01110010";
                when "1100100011" =>  -- D19.3
                    data_out_aux <= "01110011";
                when "0010110011" =>  -- D20.3
                    data_out_aux <= "01110100";
                when "1010100011" =>  -- D21.3
                    data_out_aux <= "01110101";
                when "0110100011" =>  -- D22.3
                    data_out_aux <= "01110110";
                when "0001011100" =>  -- D23.3
                    data_out_aux <= "01110111";
                when "0011001100" =>  -- D24.3
                    data_out_aux <= "01111000";
                when "1001100011" =>  -- D25.3
                    data_out_aux <= "01111001";
                when "0101100011" =>  -- D26.3
                    data_out_aux <= "01111010";
                when "0010011100" =>  -- D27.3
                    data_out_aux <= "01111011";
                when "0011100011" =>  -- D28.3
                    data_out_aux <= "01111100";
                when "0100011100" =>  -- D29.3
                    data_out_aux <= "01111101";
                when "1000011100" =>  -- D30.3
                    data_out_aux <= "01111110";
                when "0101001100" =>  -- D31.3
                    data_out_aux <= "01111111";
                when "0110001101" =>  -- D0.4
                    data_out_aux <= "10000000";
                when "1000101101" =>  -- D1.4
                    data_out_aux <= "10000001";
                when "0100101101" =>  -- D2.4
                    data_out_aux <= "10000010";
                when "1100010010" =>  -- D3.4
                    data_out_aux <= "10000011";
                when "0010101101" =>  -- D4.4
                    data_out_aux <= "10000100";
                when "1010010010" =>  -- D5.4
                    data_out_aux <= "10000101";
                when "0110010010" =>  -- D6.4
                    data_out_aux <= "10000110";
                when "0001110010" =>  -- D7.4
                    data_out_aux <= "10000111";
                when "0001101101" =>  -- D8.4
                    data_out_aux <= "10001000";
                when "1001010010" =>  -- D9.4
                    data_out_aux <= "10001001";
                when "0101010010" =>  -- D10.4
                    data_out_aux <= "10001010";
                when "1101000010" =>  -- D11.4
                    data_out_aux <= "10001011";
                when "0011010010" =>  -- D12.4
                    data_out_aux <= "10001100";
                when "1011000010" =>  -- D13.4
                    data_out_aux <= "10001101";
                when "0111000010" =>  -- D14.4
                    data_out_aux <= "10001110";
                when "1010001101" =>  -- D15.4
                    data_out_aux <= "10001111";
                when "1001001101" =>  -- D16.4
                    data_out_aux <= "10010000";
                when "1000110010" =>  -- D17.4
                    data_out_aux <= "10010001";
                when "0100110010" =>  -- D18.4
                    data_out_aux <= "10010010";
                when "1100100010" =>  -- D19.4
                    data_out_aux <= "10010011";
                when "0010110010" =>  -- D20.4
                    data_out_aux <= "10010100";
                when "1010100010" =>  -- D21.4
                    data_out_aux <= "10010101";
                when "0110100010" =>  -- D22.4
                    data_out_aux <= "10010110";
                when "0001011101" =>  -- D23.4
                    data_out_aux <= "10010111";
                when "0011001101" =>  -- D24.4
                    data_out_aux <= "10011000";
                when "1001100010" =>  -- D25.4
                    data_out_aux <= "10011001";
                when "0101100010" =>  -- D26.4
                    data_out_aux <= "10011010";
                when "0010011101" =>  -- D27.4
                    data_out_aux <= "10011011";
                when "0011100010" =>  -- D28.4
                    data_out_aux <= "10011100";
                when "0100011101" =>  -- D29.4
                    data_out_aux <= "10011101";
                when "1000011101" =>  -- D30.4
                    data_out_aux <= "10011110";
                when "0101001101" =>  -- D31.4
                    data_out_aux <= "10011111";
                when "0110001010" =>  -- D0.5
                    data_out_aux <= "10100000";
                when "1000101010" =>  -- D1.5
                    data_out_aux <= "10100001";
                when "0100101010" =>  -- D2.5
                    data_out_aux <= "10100010";
                when "1100011010" =>  -- D3.5
                    data_out_aux <= "10100011";
                when "0010101010" =>  -- D4.5
                    data_out_aux <= "10100100";
                when "1010011010" =>  -- D5.5
                    data_out_aux <= "10100101";
                when "0110011010" =>  -- D6.5
                    data_out_aux <= "10100110";
                when "0001111010" =>  -- D7.5
                    data_out_aux <= "10100111";
                when "0001101010" =>  -- D8.5
                    data_out_aux <= "10101000";
                when "1001011010" =>  -- D9.5
                    data_out_aux <= "10101001";
                when "0101011010" =>  -- D10.5
                    data_out_aux <= "10101010";
                when "1101001010" =>  -- D11.5
                    data_out_aux <= "10101011";
                when "0011011010" =>  -- D12.5
                    data_out_aux <= "10101100";
                when "1011001010" =>  -- D13.5
                    data_out_aux <= "10101101";
                when "0111001010" =>  -- D14.5
                    data_out_aux <= "10101110";
                when "1010001010" =>  -- D15.5
                    data_out_aux <= "10101111";
                when "1001001010" =>  -- D16.5
                    data_out_aux <= "10110000";
                when "1000111010" =>  -- D17.5
                    data_out_aux <= "10110001";
                when "0100111010" =>  -- D18.5
                    data_out_aux <= "10110010";
                when "1100101010" =>  -- D19.5
                    data_out_aux <= "10110011";
                when "0010111010" =>  -- D20.5
                    data_out_aux <= "10110100";
                when "1010101010" =>  -- D21.5
                    data_out_aux <= "10110101";
                when "0110101010" =>  -- D22.5
                    data_out_aux <= "10110110";
                when "0001011010" =>  -- D23.5
                    data_out_aux <= "10110111";
                when "0011001010" =>  -- D24.5
                    data_out_aux <= "10111000";
                when "1001101010" =>  -- D25.5
                    data_out_aux <= "10111001";
                when "0101101010" =>  -- D26.5
                    data_out_aux <= "10111010";
                when "0010011010" =>  -- D27.5
                    data_out_aux <= "10111011";
                when "0011101010" =>  -- D28.5
                    data_out_aux <= "10111100";
                when "0100011010" =>  -- D29.5
                    data_out_aux <= "10111101";
                when "1000011010" =>  -- D30.5
                    data_out_aux <= "10111110";
                when "0101001010" =>  -- D31.5
                    data_out_aux <= "10111111";
                when "0110000110" =>  -- D0.6
                    data_out_aux <= "11000000";
                when "1000100110" =>  -- D1.6
                    data_out_aux <= "11000001";
                when "0100100110" =>  -- D2.6
                    data_out_aux <= "11000010";
                when "1100010110" =>  -- D3.6
                    data_out_aux <= "11000011";
                when "0010100110" =>  -- D4.6
                    data_out_aux <= "11000100";
                when "1010010110" =>  -- D5.6
                    data_out_aux <= "11000101";
                when "0110010110" =>  -- D6.6
                    data_out_aux <= "11000110";
                when "0001110110" =>  -- D7.6
                    data_out_aux <= "11000111";
                when "0001100110" =>  -- D8.6
                    data_out_aux <= "11001000";
                when "1001010110" =>  -- D9.6
                    data_out_aux <= "11001001";
                when "0101010110" =>  -- D10.6
                    data_out_aux <= "11001010";
                when "1101000110" =>  -- D11.6
                    data_out_aux <= "11001011";
                when "0011010110" =>  -- D12.6
                    data_out_aux <= "11001100";
                when "1011000110" =>  -- D13.6
                    data_out_aux <= "11001101";
                when "0111000110" =>  -- D14.6
                    data_out_aux <= "11001110";
                when "1010000110" =>  -- D15.6
                    data_out_aux <= "11001111";
                when "1001000110" =>  -- D16.6
                    data_out_aux <= "11010000";
                when "1000110110" =>  -- D17.6
                    data_out_aux <= "11010001";
                when "0100110110" =>  -- D18.6
                    data_out_aux <= "11010010";
                when "1100100110" =>  -- D19.6
                    data_out_aux <= "11010011";
                when "0010110110" =>  -- D20.6
                    data_out_aux <= "11010100";
                when "1010100110" =>  -- D21.6
                    data_out_aux <= "11010101";
                when "0110100110" =>  -- D22.6
                    data_out_aux <= "11010110";
                when "0001010110" =>  -- D23.6
                    data_out_aux <= "11010111";
                when "0011000110" =>  -- D24.6
                    data_out_aux <= "11011000";
                when "1001100110" =>  -- D25.6
                    data_out_aux <= "11011001";
                when "0101100110" =>  -- D26.6
                    data_out_aux <= "11011010";
                when "0010010110" =>  -- D27.6
                    data_out_aux <= "11011011";
                when "0011100110" =>  -- D28.6
                    data_out_aux <= "11011100";
                when "0100010110" =>  -- D29.6
                    data_out_aux <= "11011101";
                when "1000010110" =>  -- D30.6
                    data_out_aux <= "11011110";
                when "0101000110" =>  -- D31.6
                    data_out_aux <= "11011111";
                when "0110001110" =>  -- D0.7
                    data_out_aux <= "11100000";
                when "1000101110" =>  -- D1.7
                    data_out_aux <= "11100001";
                when "0100101110" =>  -- D2.7
                    data_out_aux <= "11100010";
                when "1100010001" =>  -- D3.7
                    data_out_aux <= "11100011";
                when "0010101110" =>  -- D4.7
                    data_out_aux <= "11100100";
                when "1010010001" =>  -- D5.7
                    data_out_aux <= "11100101";
                when "0110010001" =>  -- D6.7
                    data_out_aux <= "11100110";
                when "0001110001" =>  -- D7.7
                    data_out_aux <= "11100111";
                when "0001101110" =>  -- D8.7
                    data_out_aux <= "11101000";
                when "1001010001" =>  -- D9.7
                    data_out_aux <= "11101001";
                when "0101010001" =>  -- D10.7
                    data_out_aux <= "11101010";
                when "1101001000" =>  -- D11.7
                    data_out_aux <= "11101011";
                when "0011010001" =>  -- D12.7
                    data_out_aux <= "11101100";
                when "1011001000" =>  -- D13.7
                    data_out_aux <= "11101101";
                when "0111001000" =>  -- D14.7
                    data_out_aux <= "11101110";
                when "1010001110" =>  -- D15.7
                    data_out_aux <= "11101111";
                when "1001001110" =>  -- D16.7
                    data_out_aux <= "11110000";
                when "1000110001" =>  -- D17.7
                    data_out_aux <= "11110001";
                when "0100110001" =>  -- D18.7
                    data_out_aux <= "11110010";
                when "1100100001" =>  -- D19.7
                    data_out_aux <= "11110011";
                when "0010110001" =>  -- D20.7
                    data_out_aux <= "11110100";
                when "1010100001" =>  -- D21.7
                    data_out_aux <= "11110101";
                when "0110100001" =>  -- D22.7
                    data_out_aux <= "11110110";
                when "0001011110" =>  -- D23.7
                    data_out_aux <= "11110111";
                when "0011001110" =>  -- D24.7
                    data_out_aux <= "11111000";
                when "1001100001" =>  -- D25.7
                    data_out_aux <= "11111001";
                when "0101100001" =>  -- D26.7
                    data_out_aux <= "11111010";
                when "0010011110" =>  -- D27.7
                    data_out_aux <= "11111011";
                when "0011100001" =>  -- D28.7
                    data_out_aux <= "11111100";
                when "0100011110" =>  -- D29.7
                    data_out_aux <= "11111101";
                when "1000011110" =>  -- D30.7
                    data_out_aux <= "11111110";
                when "0101001110" =>  -- D31.7
                    data_out_aux <= "11111111";
                when others => 
                    data_out_aux <= (others=>'0');
            end case;
        end if;
    end process;
    
    
    data_out_aux_2 <= data_out_aux(4 downto 0) & data_out_aux(7 downto 5);
    
    process (clk, rst_n)
    begin
        if rst_n = '0' then
            data_out <= (others=>'0');
        elsif rising_edge(clk) then 
            data_out <= data_out_aux_2;
        end if;
    end process;

end arch_decoder_8b_10b;
